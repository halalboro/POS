/**
 * This file is part of the Coyote <https://github.com/fpgasystems/Coyote>
 *
 * MIT Licence
 * Copyright (c) 2021-2025, Systems Group, ETH Zurich
 * All rights reserved.
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:

 * The above copyright notice and this permission notice shall be included in all
 * copies or substantial portions of the Software.

 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
 * SOFTWARE.
 */

`timescale 1ns / 1ps

import lynxTypes::*;

`include "axi_macros.svh"
`include "lynx_macros.svh"

/**
 * @brief   Top level MMU for a single vFPGA with Memory Gateway
 *
 * Top level of a single vFPGA TLB with access control, feeds into the top level arbitration.
 *
 *  @param ID_REG       Number of associated vFPGA
 *  @param N_ENDPOINTS  Number of memory endpoints for access control
 */
module mmu_region_top #(
	parameter integer 					ID_REG = 0,
	parameter integer                   N_ENDPOINTS = 1	
) (
	// AXI tlb control and writeback
    AXI4L.s   							s_axi_ctrl_sTlb,
    AXI4L.s   							s_axi_ctrl_lTlb,

    // Control interface for memory endpoints (99 bits per endpoint)
    input logic [(99*N_ENDPOINTS)-1:0] ep_ctrl,

	// Requests user
	metaIntf.s 						    s_bpss_rd_sq,
	metaIntf.s						    s_bpss_wr_sq,

`ifdef EN_STRM
	// Stream DMAs
    dmaIntf.m                           m_rd_HDMA,
    dmaIntf.m                           m_wr_HDMA,
    metaIntf.m                          m_rd_host_done,
    metaIntf.m                          m_wr_host_done,

`ifndef EN_CRED_LOCAL
    input  logic                        rxfer_host,
    input  logic                        wxfer_host,
`endif
`endif

`ifdef EN_MEM
    // Card DMAs
    dmaIntf.m                           m_rd_DDMA [N_CARD_AXI],
    dmaIntf.m                           m_wr_DDMA [N_CARD_AXI],
    metaIntf.m                          m_rd_card_done,
    metaIntf.m                          m_wr_card_done,

`ifndef EN_CRED_LOCAL
    input  logic                        rxfer_card [N_CARD_AXI],
    input  logic                        wxfer_card [N_CARD_AXI],
`endif
`endif

    // TLB page faults (from TLB FSMs)
    metaIntf.m                          m_rd_pfault_irq,
    output logic [LEN_BITS-1:0]         m_rd_pfault_rng,
    metaIntf.s                          s_rd_pfault_ctrl,
    metaIntf.m                          m_wr_pfault_irq,
    output logic [LEN_BITS-1:0]         m_wr_pfault_rng,
    metaIntf.s                          s_wr_pfault_ctrl,

    // TLB invalidation
    metaIntf.s                          s_rd_invldt_ctrl,
    metaIntf.m                          m_rd_invldt_irq,
    metaIntf.s                          s_wr_invldt_ctrl,
    metaIntf.m                          m_wr_invldt_irq,
    
    input logic        					aclk,    
	input logic    						aresetn
);

// -- Decl -----------------------------------------------------------------------------------
// -------------------------------------------------------------------------------------------
localparam integer PG_L_SIZE = 1 << PG_L_BITS;
localparam integer PG_S_SIZE = 1 << PG_S_BITS;
localparam integer HASH_L_BITS = TLB_L_ORDER;
localparam integer HASH_S_BITS = TLB_S_ORDER;
localparam integer PHY_L_BITS = PADDR_BITS - PG_L_BITS;
localparam integer PHY_S_BITS = PADDR_BITS - PG_S_BITS;
localparam integer TAG_L_BITS = VADDR_BITS - HASH_L_BITS - PG_L_BITS;
localparam integer TAG_S_BITS = VADDR_BITS - HASH_S_BITS - PG_S_BITS;
localparam integer TLB_L_DATA_BITS = TAG_L_BITS + PID_BITS + 2 + PHY_L_BITS + HPID_BITS;
localparam integer TLB_S_DATA_BITS = TAG_S_BITS + PID_BITS + 2 + PHY_S_BITS + HPID_BITS;

// Tlb interfaces
tlbIntf #(.TLB_INTF_DATA_BITS(TLB_L_DATA_BITS)) rd_lTlb ();
tlbIntf #(.TLB_INTF_DATA_BITS(TLB_S_DATA_BITS)) rd_sTlb ();
tlbIntf #(.TLB_INTF_DATA_BITS(TLB_L_DATA_BITS)) wr_lTlb ();
tlbIntf #(.TLB_INTF_DATA_BITS(TLB_S_DATA_BITS)) wr_sTlb ();
tlbIntf #(.TLB_INTF_DATA_BITS(TLB_L_DATA_BITS)) lTlb ();
tlbIntf #(.TLB_INTF_DATA_BITS(TLB_S_DATA_BITS)) sTlb ();

AXI4S #(.AXI4S_DATA_BITS(AXI_TLB_BITS)) axis_lTlb ();
AXI4S #(.AXI4S_DATA_BITS(AXI_TLB_BITS)) axis_sTlb ();

// Request interfaces - only authorized requests from memory gateway
metaIntf #(.STYPE(req_t)) rd_req ();
metaIntf #(.STYPE(req_t)) wr_req ();

// `META_ASSIGN(s_bpss_rd_sq, rd_req)
// `META_ASSIGN(s_bpss_wr_sq, wr_req)

// ----------------------------------------------------------------------------------------
// Memory Gateway - Filters and only passes authorized requests
// ----------------------------------------------------------------------------------------
gate_mem #(
    .N_ENDPOINTS(N_ENDPOINTS)
) inst_gate_mem (
    .aclk(aclk),
    .aresetn(aresetn),
    .ep_ctrl(ep_ctrl),

    // Original user requests
    .s_rd_req(s_bpss_rd_sq),
    .s_wr_req(s_bpss_wr_sq),

    // Only authorized requests pass through to TLB FSMs
    .m_rd_req(rd_req),
    .m_wr_req(wr_req)
);

// create_ip -name ila -vendor xilinx.com -library ip -version 6.2 -module_name ila_mem_gateway
// set_property -dict [list \
//     CONFIG.C_NUM_OF_PROBES {14} \
//     CONFIG.C_PROBE0_WIDTH {1} \
//     CONFIG.C_PROBE1_WIDTH {2} \
//     CONFIG.C_PROBE2_WIDTH {64} \
//     CONFIG.C_PROBE3_WIDTH {64} \
//     CONFIG.C_PROBE4_WIDTH {64} \
//     CONFIG.C_PROBE5_WIDTH {28} \
//     CONFIG.C_PROBE6_WIDTH {64} \
//     CONFIG.C_PROBE7_WIDTH {28} \
//     CONFIG.C_PROBE8_WIDTH {1} \
//     CONFIG.C_PROBE9_WIDTH {1} \
//     CONFIG.C_PROBE10_WIDTH {1} \
//     CONFIG.C_PROBE11_WIDTH {1} \
//     CONFIG.C_PROBE12_WIDTH {1} \
//     CONFIG.C_PROBE13_WIDTH {1} \
//     CONFIG.C_EN_STRG_QUAL {1} \
//     CONFIG.ALL_PROBE_SAME_MU_CNT {2} \
// ] [get_ips ila_mem_gateway]

ila_mem_gate_signal inst_ila_mem_gate_signal (
    .clk(aclk),
    .probe0(ep_ctrl_data)
);

ila_mem_region_top_req_t inst_rd_req_ila (
    .clk(aclk),
    .probe0(s_bpss_rd_sq.data.opcode),
    .probe1(s_bpss_rd_sq.data.strm),
    .probe2(s_bpss_rd_sq.data.mode),
    .probe3(s_bpss_rd_sq.data.rdma),
    .probe4(s_bpss_rd_sq.data.remote),
    .probe5(s_bpss_rd_sq.data.vfid),
    .probe6(s_bpss_rd_sq.data.pid),
    .probe7(s_bpss_rd_sq.data.dest),
    .probe8(s_bpss_rd_sq.data.last),
    .probe9(s_bpss_rd_sq.data.vaddr),
    .probe10(s_bpss_rd_sq.data.len),
    .probe11(s_bpss_rd_sq.data.actv),
    .probe12(s_bpss_rd_sq.data.host),
    .probe13(s_bpss_rd_sq.data.offs),
    .probe14(s_bpss_rd_sq.valid),
    .probe15(s_bpss_rd_sq.ready),
    .probe16(rd_req.data.opcode),
    .probe17(rd_req.data.strm),
    .probe18(rd_req.data.mode),
    .probe19(rd_req.data.rdma),
    .probe20(rd_req.data.remote),
    .probe21(rd_req.data.vfid),
    .probe22(rd_req.data.pid),
    .probe23(rd_req.data.dest),
    .probe24(rd_req.data.last),
    .probe25(rd_req.data.vaddr),
    .probe26(rd_req.data.len),
    .probe27(rd_req.data.actv),
    .probe28(rd_req.data.host),
    .probe29(rd_req.data.offs),
    .probe30(rd_req.valid),
    .probe31(rd_req.ready)
);

// ila_mem_region_top_req_t inst_bpss_rd_req_ila (
//     .clk(aclk),
//     .probe0(s_bpss_rd_sq.data.opcode),
//     .probe1(s_bpss_rd_sq.data.strm),
//     .probe2(s_bpss_rd_sq.data.mode),
//     .probe3(s_bpss_rd_sq.data.rdma),
//     .probe4(s_bpss_rd_sq.data.remote),
//     .probe5(s_bpss_rd_sq.data.vfid),
//     .probe6(s_bpss_rd_sq.data.pid),
//     .probe7(s_bpss_rd_sq.data.dest),
//     .probe8(s_bpss_rd_sq.data.last),
//     .probe9(s_bpss_rd_sq.data.vaddr),
//     .probe10(s_bpss_rd_sq.data.len),
//     .probe11(s_bpss_rd_sq.data.actv),
//     .probe12(s_bpss_rd_sq.data.host),
//     .probe13(s_bpss_rd_sq.data.offs),
//     .probe14(s_bpss_rd_sq.valid),
//     .probe15(s_bpss_rd_sq.ready)
// );

// ila_mem_region_top_req_t inst_rd_req_ila (
//     .clk(aclk),
//     .probe0(rd_req.data.opcode),
//     .probe1(rd_req.data.strm),
//     .probe2(rd_req.data.mode),
//     .probe3(rd_req.data.rdma),
//     .probe4(rd_req.data.remote),
//     .probe5(rd_req.data.vfid),
//     .probe6(rd_req.data.pid),
//     .probe7(rd_req.data.dest),
//     .probe8(rd_req.data.last),
//     .probe9(rd_req.data.vaddr),
//     .probe10(rd_req.data.len),
//     .probe11(rd_req.data.actv),
//     .probe12(rd_req.data.host),
//     .probe13(rd_req.data.offs),
//     .probe14(rd_req.valid),
//     .probe15(rd_req.ready)
// );

// ----------------------------------------------------------------------------------------
// Mutex 
// ----------------------------------------------------------------------------------------
logic [1:0] mutex;
logic rd_lock, wr_lock;
logic rd_unlock, wr_unlock;

always_ff @(posedge aclk) begin
	if(aresetn == 1'b0) begin
		mutex <= 2'b01;
	end else begin
		if(mutex[0] == 1'b1) begin // free
			if(rd_lock)
				mutex <= 2'b00;
			else if(wr_lock)
				mutex <= 2'b10;
		end
		else begin // locked
			if((mutex[1] == 1'b0) && rd_unlock)
				mutex <= 2'b01;
			else if (wr_unlock)
				mutex <= 2'b11;
		end
	end
end

// ----------------------------------------------------------------------------------------
// TLB
// ---------------------------------------------------------------------------------------- 
assign rd_lTlb.data = lTlb.data;
assign wr_lTlb.data = lTlb.data;
assign rd_sTlb.data = sTlb.data;
assign wr_sTlb.data = sTlb.data;
assign rd_lTlb.hit  = lTlb.hit;
assign wr_lTlb.hit  = lTlb.hit;
assign rd_sTlb.hit  = sTlb.hit;
assign wr_sTlb.hit  = sTlb.hit;

assign lTlb.addr  = mutex[1] ? wr_lTlb.addr : rd_lTlb.addr;
assign sTlb.addr  = mutex[1] ? wr_sTlb.addr : rd_sTlb.addr;
assign lTlb.pid   = mutex[1] ? wr_lTlb.pid : rd_lTlb.pid;
assign sTlb.pid   = mutex[1] ? wr_sTlb.pid : rd_sTlb.pid;
assign lTlb.strm  = mutex[1] ? wr_lTlb.strm : rd_lTlb.strm;
assign sTlb.strm  = mutex[1] ? wr_sTlb.strm : rd_sTlb.strm;
assign lTlb.wr    = mutex[1] ? wr_lTlb.wr : rd_lTlb.wr;
assign sTlb.wr    = mutex[1] ? wr_sTlb.wr : rd_sTlb.wr;
assign lTlb.valid = mutex[1] ? wr_lTlb.valid : rd_lTlb.valid;
assign sTlb.valid = mutex[1] ? wr_sTlb.valid : rd_sTlb.valid;

// TLBs
tlb_controller #(
    .TLB_ORDER(TLB_L_ORDER),
    .PG_BITS(PG_L_BITS),
    .N_ASSOC(N_L_ASSOC),
    .DBG_L(1),
    .ID_REG(ID_REG)
) inst_lTlb (
    .aclk(aclk),
    .aresetn(aresetn),
    .s_axis(axis_lTlb),
    .TLB(lTlb)
);

tlb_controller #(
    .TLB_ORDER(TLB_S_ORDER),
    .PG_BITS(PG_S_BITS),
    .N_ASSOC(N_S_ASSOC),
    .DBG_S(1),
    .ID_REG(ID_REG)
) inst_sTlb (
    .aclk(aclk),
    .aresetn(aresetn),
    .s_axis(axis_sTlb),
    .TLB(sTlb)
);

// TLB slaves
tlb_slave_axil #(
    .TLB_ORDER(TLB_L_ORDER),
    .PG_BITS(PG_L_BITS),
    .N_ASSOC(N_L_ASSOC)
) inst_lTlb_slv_0 (
    .aclk(aclk),
    .aresetn(aresetn),
    .s_axi_ctrl(s_axi_ctrl_lTlb),
    .m_axis(axis_lTlb)
);

tlb_slave_axil #(
    .TLB_ORDER(TLB_S_ORDER),
    .PG_BITS(PG_S_BITS),
    .N_ASSOC(N_S_ASSOC)
) inst_sTlb_slv_0 (
    .aclk(aclk),
    .aresetn(aresetn),
    .s_axi_ctrl(s_axi_ctrl_sTlb),
    .m_axis(axis_sTlb)
);

// ----------------------------------------------------------------------------------------
// FSM
// ----------------------------------------------------------------------------------------
`ifdef EN_STRM
    // FSM
    dmaIntf rd_HDMA_fsm ();
    dmaIntf wr_HDMA_fsm ();
    
    // Queue
    dmaIntf rd_HDMA_fsm_q ();
    dmaIntf wr_HDMA_fsm_q ();

    // Parsing
    dmaIntf rd_HDMA_parsed ();
    dmaIntf wr_HDMA_parsed ();

    // Credits
    dmaIntf rd_HDMA_cred ();
    dmaIntf wr_HDMA_cred ();
`endif

`ifdef EN_MEM
    // FSM
    dmaIntf rd_DDMA_fsm [N_CARD_AXI] ();
    dmaIntf wr_DDMA_fsm [N_CARD_AXI] ();

    // Queue
    dmaIntf rd_DDMA_fsm_q [N_CARD_AXI] ();
    dmaIntf wr_DDMA_fsm_q [N_CARD_AXI] ();

    // Parsing
    dmaIntf rd_DDMA_parsed [N_CARD_AXI] ();
    dmaIntf wr_DDMA_parsed [N_CARD_AXI] ();

    // Credits
    dmaIntf rd_DDMA_cred [N_CARD_AXI] ();
    dmaIntf wr_DDMA_cred [N_CARD_AXI] ();
`endif

// TLB rd FSM - receives only authorized requests
tlb_fsm #(
    .ID_REG(ID_REG),
    .RDWR(0)
) inst_fsm_rd (
    .aclk(aclk),
    .aresetn(aresetn),
    .lTlb(rd_lTlb),
    .sTlb(rd_sTlb),
`ifdef EN_STRM
    .m_host_done(m_rd_host_done),
    .m_HDMA(rd_HDMA_fsm),
`endif
`ifdef EN_MEM
    .m_card_done(m_rd_card_done),
    .m_DDMA(rd_DDMA_fsm),
`endif
    .s_req(rd_req),  // Only authorized requests from memory gateway

    .m_pfault(m_rd_pfault_irq),
    .m_pfault_rng(m_rd_pfault_rng),
    .s_pfault(s_rd_pfault_ctrl),

    .s_invldt(s_rd_invldt_ctrl),
    .m_invldt(m_rd_invldt_irq),

    .lock(rd_lock),
	.unlock(rd_unlock),
	.mutex(mutex)
);

// TLB wr FSM - receives only authorized requests
tlb_fsm #(
    .ID_REG(ID_REG),
    .RDWR(1)
) inst_fsm_wr (
    .aclk(aclk),
    .aresetn(aresetn),
    .lTlb(wr_lTlb),
    .sTlb(wr_sTlb),
`ifdef EN_STRM
    .m_host_done(m_wr_host_done),
    .m_HDMA(wr_HDMA_fsm),
`endif
`ifdef EN_MEM
    .m_card_done(m_wr_card_done),
    .m_DDMA(wr_DDMA_fsm),
`endif
    .s_req(wr_req),  // Only authorized requests from memory gateway

    .m_pfault(m_wr_pfault_irq),
    .m_pfault_rng(m_wr_pfault_rng),
    .s_pfault(s_wr_pfault_ctrl),

    .s_invldt(s_wr_invldt_ctrl),
    .m_invldt(m_wr_invldt_irq),

    .lock(wr_lock),
	.unlock(wr_unlock),
	.mutex(mutex)
);

// ----------------------------------------------------------------------------------------
// Queueing stage
// ----------------------------------------------------------------------------------------
`ifdef EN_STRM
    // HDMA
    dma_req_queue inst_rd_q_fsm_hdma (.aclk(aclk), .aresetn(aresetn), .s_req(rd_HDMA_fsm), .m_req(rd_HDMA_fsm_q));
    dma_req_queue inst_wr_q_fsm_hdma (.aclk(aclk), .aresetn(aresetn), .s_req(wr_HDMA_fsm), .m_req(wr_HDMA_fsm_q));

    // Parsing 
`ifndef EN_CRED_LOCAL
    dma_parser inst_rd_parser (.aclk(aclk), .aresetn(aresetn), .s_req(rd_HDMA_fsm_q), .m_req(rd_HDMA_parsed));
    dma_parser inst_wr_parser (.aclk(aclk), .aresetn(aresetn), .s_req(wr_HDMA_fsm_q), .m_req(wr_HDMA_parsed));
`else
    `DMA_REQ_ASSIGN(rd_HDMA_fsm_q, rd_HDMA_parsed)
    `DMA_REQ_ASSIGN(wr_HDMA_fsm_q, wr_HDMA_parsed)
`endif
`endif

`ifdef EN_MEM
    for(genvar i = 0; i < N_CARD_AXI; i++) begin
        // DDMA
        dma_req_queue inst_rd_q_fsm_ddma (.aclk(aclk), .aresetn(aresetn), .s_req(rd_DDMA_fsm[i]), .m_req(rd_DDMA_fsm_q[i]));
        dma_req_queue inst_wr_q_fsm_ddma (.aclk(aclk), .aresetn(aresetn), .s_req(wr_DDMA_fsm[i]), .m_req(wr_DDMA_fsm_q[i]));
    end

    // Parsing 
`ifndef EN_CRED_LOCAL
    for(genvar i = 0; i < N_CARD_AXI; i++) begin
        dma_parser inst_rd_parser (.aclk(aclk), .aresetn(aresetn), .s_req(rd_DDMA_fsm_q[i]), .m_req(rd_DDMA_parsed[i]));
        dma_parser inst_wr_parser (.aclk(aclk), .aresetn(aresetn), .s_req(wr_DDMA_fsm_q[i]), .m_req(wr_DDMA_parsed[i]));
    end
`else
    for(genvar i = 0; i < N_CARD_AXI; i++) begin
        `DMA_REQ_ASSIGN(rd_DDMA_fsm_q[i], rd_DDMA_parsed[i])
        `DMA_REQ_ASSIGN(wr_DDMA_fsm_q[i], wr_DDMA_parsed[i])
    end
`endif
`endif

// ----------------------------------------------------------------------------------------
// Credits and output
// ----------------------------------------------------------------------------------------
`ifndef EN_CRED_LOCAL

`ifdef EN_STRM
    // HDMA
    mmu_credits_rd #(.ID_REG(ID_REG)) inst_rd_cred_hdma (.aclk(aclk), .aresetn(aresetn), .s_req(rd_HDMA_parsed), .m_req(rd_HDMA_cred), .rxfer(rxfer_host));
    mmu_credits_wr #(.ID_REG(ID_REG)) inst_wr_cred_hdma (.aclk(aclk), .aresetn(aresetn), .s_req(wr_HDMA_parsed), .m_req(wr_HDMA_cred), .wxfer(wxfer_host));

    // Queueing
    dma_req_queue inst_rd_q_cred_hdma (.aclk(aclk), .aresetn(aresetn), .s_req(rd_HDMA_cred), .m_req(m_rd_HDMA));
    dma_req_queue inst_wr_q_cred_hdma (.aclk(aclk), .aresetn(aresetn), .s_req(wr_HDMA_cred), .m_req(m_wr_HDMA));
`endif

`ifdef EN_MEM
    for(genvar i = 0; i < N_CARD_AXI; i++) begin
        // DDMA
        mmu_credits_rd #(.ID_REG(ID_REG)) inst_rd_cred_ddma (.aclk(aclk), .aresetn(aresetn), .s_req(rd_DDMA_parsed[i]), .m_req(rd_DDMA_cred[i]), .rxfer(rxfer_card[i]));
        mmu_credits_wr #(.ID_REG(ID_REG)) inst_wr_cred_ddma (.aclk(aclk), .aresetn(aresetn), .s_req(wr_DDMA_parsed[i]), .m_req(wr_DDMA_cred[i]), .wxfer(wxfer_card[i]));

        // Queueing
        dma_req_queue inst_rd_q_cred_ddma (.aclk(aclk), .aresetn(aresetn), .s_req(rd_DDMA_cred[i]), .m_req(m_rd_DDMA[i]));
        dma_req_queue inst_wr_q_cred_ddma (.aclk(aclk), .aresetn(aresetn), .s_req(wr_DDMA_cred[i]), .m_req(m_wr_DDMA[i]));
    end
`endif

`else

`ifdef EN_STRM
    `DMA_REQ_ASSIGN(rd_HDMA_parsed, m_rd_HDMA)
    `DMA_REQ_ASSIGN(wr_HDMA_parsed, m_wr_HDMA)
`endif

`ifdef EN_MEM
    for(genvar i = 0; i < N_CARD_AXI; i++) begin
        `DMA_REQ_ASSIGN(rd_DDMA_parsed[i], m_rd_DDMA[i])
        `DMA_REQ_ASSIGN(wr_DDMA_parsed[i], m_wr_DDMA[i])
    end
`endif

`endif

/////////////////////////////////////////////////////////////////////////////
// DEBUG
/////////////////////////////////////////////////////////////////////////////
`ifdef DBG_MMU_REGION_TOP

`endif

endmodule // mmu_region_top